`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:47:43 11/13/2014 
// Design Name: 
// Module Name:    sub_RGB 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module sub_RGB(
    input clk,
	 input ce,
    input [9:0] red,
    input [9:0] green,
    input [9:0] blue,
	 input [9:0] blue;
	 output [9:0] value,
	 output [1:0] index
    );


endmodule
