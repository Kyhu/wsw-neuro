-- Tomasz Kryjak
-- AGH Krakow

			  
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity switchModel_pbas_rgbs_19 is
	generic (
			PIXEL_W : in natural := 8;
			DIST_W  : in natural := 8;
			POS_W    : in natural := 6;
			RT_W    : in natural := 16;
			BG_MODEL_SC_W    : in natural := 336;
			BG_MODEL_ALL_W : in natural := 362
			);
    Port ( CLK : in STD_LOGIC;
			  RST : in STD_LOGIC;
			  CE : in STD_LOGIC;
			  SWITCH : in STD_LOGIC;
			  IS_CENTRAL : in STD_LOGIC;
			  TOSWITCH : in STD_LOGIC_VECTOR(7 downto 0);
           BG_MODEL_IN : in  STD_LOGIC_VECTOR (BG_MODEL_ALL_W -1 downto 0);

			  BG_MODEL_OUT : out  STD_LOGIC_VECTOR (BG_MODEL_ALL_W -1 downto 0)
			  );
end switchModel_pbas_rgbs_19;
architecture Behavioral of switchModel_pbas_rgbs_19 is
begin

	 process (CLK) is
	 begin
		 if (rising_edge(CLK) ) then
			 if ( CE = '1' ) then
				 if ( RST = '1') then
					 BG_MODEL_OUT <= (others => '0');
				 else
					 if ( SWITCH = '1' ) then

						 BG_MODEL_OUT(BG_MODEL_ALL_W -1  downto BG_MODEL_SC_W-2*RT_W) <= BG_MODEL_IN(BG_MODEL_ALL_W -1  downto BG_MODEL_SC_W-2*RT_W); 
-- UPDATE THE MIN VALUE 
						 if ( IS_CENTRAL = '1') then
							 case  BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W + POS_W -1  downto BG_MODEL_SC_W + PIXEL_W + DIST_W) is -- pos 
								 when "000000" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "000001" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "000010" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "000011" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "000100" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "000101" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "000110" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "000111" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "001000" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "001001" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "001010" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "001011" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "001100" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "001101" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "001110" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "001111" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "010000" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "010001" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(303 downto 296);
								 when "010010" => 
									 BG_MODEL_OUT(15 downto 8) <= BG_MODEL_IN(15 downto 8);
									 BG_MODEL_OUT(31 downto 24) <= BG_MODEL_IN(31 downto 24);
									 BG_MODEL_OUT(47 downto 40) <= BG_MODEL_IN(47 downto 40);
									 BG_MODEL_OUT(63 downto 56) <= BG_MODEL_IN(63 downto 56);
									 BG_MODEL_OUT(79 downto 72) <= BG_MODEL_IN(79 downto 72);
									 BG_MODEL_OUT(95 downto 88) <= BG_MODEL_IN(95 downto 88);
									 BG_MODEL_OUT(111 downto 104) <= BG_MODEL_IN(111 downto 104);
									 BG_MODEL_OUT(127 downto 120) <= BG_MODEL_IN(127 downto 120);
									 BG_MODEL_OUT(143 downto 136) <= BG_MODEL_IN(143 downto 136);
									 BG_MODEL_OUT(159 downto 152) <= BG_MODEL_IN(159 downto 152);
									 BG_MODEL_OUT(175 downto 168) <= BG_MODEL_IN(175 downto 168);
									 BG_MODEL_OUT(191 downto 184) <= BG_MODEL_IN(191 downto 184);
									 BG_MODEL_OUT(207 downto 200) <= BG_MODEL_IN(207 downto 200);
									 BG_MODEL_OUT(223 downto 216) <= BG_MODEL_IN(223 downto 216);
									 BG_MODEL_OUT(239 downto 232) <= BG_MODEL_IN(239 downto 232);
									 BG_MODEL_OUT(255 downto 248) <= BG_MODEL_IN(255 downto 248);
									 BG_MODEL_OUT(271 downto 264) <= BG_MODEL_IN(271 downto 264);
									 BG_MODEL_OUT(287 downto 280) <= BG_MODEL_IN(287 downto 280);
									 BG_MODEL_OUT(303 downto 296) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W + DIST_W -1  downto BG_MODEL_SC_W + PIXEL_W); -- minimum distance value
								 when others =>
									 BG_MODEL_OUT <= ( others => '0');
							 end case;
						 end if; 


-- UPDATE THE MODEL 
						 case  TOSWITCH  is 
							 when "00000000" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00000001" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00000010" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00000011" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00000100" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00000101" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00000110" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00000111" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00001000" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00001001" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00001010" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00001011" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00001100" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00001101" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00001110" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00001111" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00010000" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00010001" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(295 downto 288);
							 when "00010010" => 
								 BG_MODEL_OUT(7 downto 0) <= BG_MODEL_IN(7 downto 0);
								 BG_MODEL_OUT(23 downto 16) <= BG_MODEL_IN(23 downto 16);
								 BG_MODEL_OUT(39 downto 32) <= BG_MODEL_IN(39 downto 32);
								 BG_MODEL_OUT(55 downto 48) <= BG_MODEL_IN(55 downto 48);
								 BG_MODEL_OUT(71 downto 64) <= BG_MODEL_IN(71 downto 64);
								 BG_MODEL_OUT(87 downto 80) <= BG_MODEL_IN(87 downto 80);
								 BG_MODEL_OUT(103 downto 96) <= BG_MODEL_IN(103 downto 96);
								 BG_MODEL_OUT(119 downto 112) <= BG_MODEL_IN(119 downto 112);
								 BG_MODEL_OUT(135 downto 128) <= BG_MODEL_IN(135 downto 128);
								 BG_MODEL_OUT(151 downto 144) <= BG_MODEL_IN(151 downto 144);
								 BG_MODEL_OUT(167 downto 160) <= BG_MODEL_IN(167 downto 160);
								 BG_MODEL_OUT(183 downto 176) <= BG_MODEL_IN(183 downto 176);
								 BG_MODEL_OUT(199 downto 192) <= BG_MODEL_IN(199 downto 192);
								 BG_MODEL_OUT(215 downto 208) <= BG_MODEL_IN(215 downto 208);
								 BG_MODEL_OUT(231 downto 224) <= BG_MODEL_IN(231 downto 224);
								 BG_MODEL_OUT(247 downto 240) <= BG_MODEL_IN(247 downto 240);
								 BG_MODEL_OUT(263 downto 256) <= BG_MODEL_IN(263 downto 256);
								 BG_MODEL_OUT(279 downto 272) <= BG_MODEL_IN(279 downto 272);
								 BG_MODEL_OUT(295 downto 288) <= BG_MODEL_IN(BG_MODEL_SC_W + PIXEL_W -1  downto BG_MODEL_SC_W); -- PIXEL;
							 when others =>
								 BG_MODEL_OUT <= ( others => '0');
						 end case;
					 else
						 BG_MODEL_OUT <= BG_MODEL_IN;
					 end if;
				 end if;		
			 end if;	
		 end if;	
	 end process;


end Behavioral;
